---------------------------------------------------------------------
--
-- Built with PASM version 1.3
-- File name: myco_mem.vhd
-- 8-7-2023 20:20:49
-- 
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity myco_mem is
port (
    clock        : in std_logic;
    clock_enable : in std_logic;
    address      : in std_logic_vector(9 downto 0);
    data_out     : out std_logic_vector(15 downto 0);
    data_in      : in std_logic_vector(15 downto 0);
    write_enable : in std_logic);
end entity;

architecture rtl of myco_mem is

    type ram_type is array (0 to 1023) of std_logic_vector(15 downto 0);
    signal ram : ram_type := (
			X"B012",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0001",X"0002",
			X"0003",X"0004",X"0221",X"1001",X"1002",X"1003",X"1004",X"1006",
			X"1007",X"A011",X"A00E",X"900D",X"100C",X"5222",X"D029",X"1005",
			X"A00E",X"0223",X"A010",X"E0A5",X"E041",X"E04F",X"0005",X"2224",
			X"B01F",X"0221",X"1005",X"E0A5",X"0225",X"2009",X"4226",X"1030",
			X"B031",X"B0AF",X"B0B2",X"B0B5",X"B0CB",X"B0CE",X"B0D1",X"B104",
			X"B130",X"B17D",X"B182",X"B185",X"B18A",X"B18F",X"B1DB",X"B1DE",
			X"B0AF",X"0009",X"A00E",X"E082",X"D04E",X"0221",X"1009",X"A00E",
			X"E05D",X"E082",X"D04E",X"0009",X"2224",X"B046",X"F000",X"0008",
			X"A00E",X"E082",X"D05C",X"0221",X"1008",X"A00E",X"E05D",X"E082",
			X"D05C",X"0008",X"2224",X"B054",X"F000",X"0009",X"100B",X"E086",
			X"4008",X"100A",X"E07C",X"000A",X"100B",X"E075",X"7005",X"0227",
			X"C06A",X"0228",X"500A",X"400B",X"100A",X"7005",X"5229",X"222A",
			X"422B",X"1073",X"000A",X"B074",X"F000",X"7005",X"5229",X"222A",
			X"1079",X"B07A",X"100A",X"F000",X"7005",X"C07F",X"F000",X"800A",
			X"100A",X"F000",X"E093",X"3224",X"C082",X"F000",X"E089",X"E089",
			X"E089",X"000B",X"200B",X"100B",X"F000",X"E090",X"E090",X"E090",
			X"700A",X"100A",X"F000",X"900D",X"600C",X"D098",X"0221",X"F000",
			X"100A",X"022C",X"A010",X"900D",X"600C",X"600A",X"D096",X"000A",
			X"600C",X"100C",X"622D",X"500A",X"F000",X"E075",X"E07C",X"000A",
			X"522E",X"1008",X"E08D",X"000A",X"522E",X"1009",X"F000",X"0005",
			X"2224",X"B02A",X"0008",X"A00E",X"B0AF",X"022F",X"2008",X"10B8",
			X"B0B9",X"A010",X"B0AF",X"0001",X"0002",X"0005",X"000A",X"0014",
			X"0032",X"0064",X"00C8",X"01F4",X"03E8",X"07D0",X"1388",X"2710",
			X"4E20",X"7530",X"EA60",X"0005",X"3008",X"B02A",X"0008",X"1001",
			X"B0AF",X"0230",X"2008",X"4226",X"10D6",X"0001",X"B0D7",X"B0AF",
			X"B0E7",X"B0E9",X"B0EB",X"B0ED",X"B0EF",X"B0F1",X"B0F3",X"B0F5",
			X"B102",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"1002",
			X"B0AF",X"1003",X"B0AF",X"1004",X"B0AF",X"A00E",X"B0AF",X"0224",
			X"B0F6",X"0222",X"B0F6",X"0231",X"B0F6",X"0232",X"100A",X"7001",
			X"C0FC",X"900E",X"400A",X"B0ED",X"000A",X"622E",X"100A",X"900E",
			X"500A",X"B0ED",X"A011",X"B0AF",X"0233",X"2008",X"4226",X"1109",
			X"900F",X"B10A",X"B0AF",X"B11A",X"B11D",X"B11F",X"B121",X"B123",
			X"B125",X"B127",X"B129",X"B12E",X"B12E",X"B0AF",X"B0AF",X"B0AF",
			X"B0AF",X"B0AF",X"0002",X"1001",X"B0AF",X"0003",X"B11B",X"0004",
			X"B11B",X"900F",X"B11B",X"5224",X"B12A",X"5222",X"B12A",X"5231",
			X"B12A",X"5232",X"D12C",X"B11B",X"0224",X"B11B",X"0221",X"B11B",
			X"0234",X"2008",X"4226",X"1135",X"0001",X"B136",X"B0AF",X"B146",
			X"B149",X"B14B",X"B14D",X"B14F",X"B163",X"B175",X"B177",X"B179",
			X"B17B",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"2224",X"1001",
			X"B0AF",X"3224",X"B147",X"2002",X"B147",X"3002",X"B147",X"0002",
			X"100B",X"E086",X"0231",X"100A",X"000B",X"200B",X"100B",X"5235",
			X"D15A",X"B15D",X"000B",X"2001",X"100B",X"000A",X"3224",X"D153",
			X"000B",X"522E",X"B147",X"0002",X"100B",X"E086",X"0231",X"100A",
			X"0001",X"2001",X"1001",X"300B",X"C16F",X"4224",X"1001",X"000A",
			X"3224",X"D167",X"0001",X"522E",X"B147",X"5002",X"B147",X"4002",
			X"B147",X"6002",X"B147",X"622E",X"B147",X"0008",X"100B",X"E086",
			X"1006",X"B0AF",X"0006",X"4008",X"B02A",X"0003",X"3224",X"C0AF",
			X"1003",X"B182",X"0004",X"3224",X"C0AF",X"1004",X"B182",X"0236",
			X"2008",X"4226",X"1193",X"B194",X"B0AF",X"B1A4",X"B1A8",X"B1AC",
			X"B1B0",X"B1B2",X"B1B4",X"B1B6",X"B1BC",X"B1BE",X"B1C0",X"B1C2",
			X"B1C8",X"B1CC",X"B1D0",X"B1D4",X"0002",X"3001",X"C1D8",X"B0AF",
			X"0001",X"3002",X"C1D8",X"B0AF",X"0001",X"3002",X"D0AF",X"B1D8",
			X"0224",X"B1B7",X"0222",X"B1B7",X"0231",X"B1B7",X"0232",X"100B",
			X"900F",X"500B",X"D1D8",X"B0AF",X"0224",X"B1C3",X"0222",X"B1C3",
			X"0231",X"B1C3",X"0232",X"100B",X"900F",X"500B",X"D0AF",X"B1D8",
			X"900D",X"5224",X"D0AF",X"B1D8",X"900D",X"5222",X"D0AF",X"B1D8",
			X"900D",X"5224",X"D1D8",X"B0AF",X"900D",X"5222",X"D1D8",X"B0AF",
			X"0005",X"2222",X"B02A",X"0005",X"1007",X"B182",X"0007",X"1005",
			X"B0AF",X"6451",X"4E80",X"C398",X"8295",X"4D80",X"C39E",X"829A",
			X"4B81",X"C394",X"8390",X"4781",X"C39A",X"8394",X"4382",X"C390",
			X"8490",X"1128",X"1828",X"3471",X"5459",X"2634",X"6954",X"5926",
			X"34FF",X"54CE",X"7133",X"22CC",X"3240",X"2271",X"54CE",X"3439",
			X"FFFF",X"86D0",X"4071",X"5423",X"CD34",X"D840",X"543B",X"FFFF",
			X"FFFF",X"4F93",X"4553",X"1911",X"2119",X"1121",X"1911",X"20B4",
			X"10E0",X"23CE",X"3223",X"CC31",X"E0FF",X"23CF",X"3223",X"CD31",
			X"E0FF",X"CC31",X"4054",X"23CE",X"32CF",X"E0CC",X"3371",X"23CC",
			X"313C",X"0000",X"0002",X"012C",X"0001",X"0031",X"B000",X"00FF",
			X"FF00",X"003F",X"01E1",X"1000",X"001E",X"0003",X"000F",X"00BB",
			X"00D7",X"0004",X"0008",X"010A",X"0136",X"0100",X"0194",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000");
begin

    process(clock)
    begin
        if rising_edge(clock) then
            if clock_enable = '1' then
                if write_enable = '1' then
                    ram(to_integer(unsigned(address))) <= data_in;
                else
                    data_out <= ram(to_integer(unsigned(address)));
                end if;
            end if;
        end if;
    end process;

end rtl;

--- End of file ---
